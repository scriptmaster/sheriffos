module main

fn main() {
	println(c'hi')
}
